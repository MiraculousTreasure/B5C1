terminal id :ssh -X Pyadav@172.16.17.6
